
netcdf mir_scld1c_organised_by_snapshot {
dimensions:
    snapshot_counter = unlimited ; // actual value is the number of snapshots in original file
    grid_point_counter = 2400 ; // or whatever the maximum number of grid points per snapshot is, always this value
    radiometric_accuracy_counter = 2; // always this value
variables:
    unsigned short grid_point_counter(snapshot_counter) ;
    unsigned int grid_point_id(snapshot_counter, grid_point_counter) ;
    float grid_point_latitude(snapshot_counter, grid_point_counter) ;
        grid_point_latitude:units = "degrees_north" ;
        grid_point_latitude:_FillValue = -999.f ;
        grid_point_latitude:valid_min = -90.f ;
        grid_point_latitude:valid_max = 90.f ;
    float grid_point_longitude(snapshot_counter, grid_point_counter) ;
        grid_point_longitude:units = "degrees_east" ;
        grid_point_longitude:_FillValue = -999.f ;
        grid_point_longitude:valid_min = -180.f ;
        grid_point_longitude:valid_max = 180.f ;
    float grid_point_altitude(snapshot_counter, grid_point_counter) ;
        grid_point_altitude:units = “m” ;
        grid_point_altitude:_FillValue = -999.f ;
    unsigned byte grid_point_mask(snapshot_counter, grid_point_counter) ;
    unsigned short bt_data_counter(snapshot_counter, grid_point_counter) ;
    unsigned short flags(snapshot_counter, grid_point_counter) ;
    unsigned float bt_value(snapshot_counter, grid_point_counter) ;
    unsigned short pixel_radiometric_accuracy(snapshot_counter, grid_point_counter) ;
    unsigned short incidence_angle(snapshot_counter, grid_point_counter) ;
    unsigned short azimuth_angle(snapshot_counter, grid_point_counter) ;
    unsigned short faraday_rotation_angle(snapshot_counter, grid_point_counter) ;
    unsigned short geometric_rotation_angle(snapshot_counter, grid_point_counter) ;
    // unsigned int snapshot_id_of_pixel(snapshot_counter, grid_point_counter) ;
    unsigned short footprint_axis_1(snapshot_counter, grid_point_counter) ;
    unsigned short footprint_axis_2(snapshot_counter, grid_point_counter) ;

    int snapshot_time_days(snapshot_counter) ;
    unsigned int snapshot_time_seconds(snapshot_counter) ;
    unsigned int snapshot_time_microseconds(snapshot_counter) ;
    unsigned int snapshot_id(snapshot_counter) ;
    unsigned long long snapshot_obet(snapshot_counter) ;    
    double x_position(snapshot_counter);
    double y_position(snapshot_counter);
    double z_position(snapshot_counter);
    double x_velocity(snapshot_counter);
    double y_velocity(snapshot_counter);
    double z_velocity(snapshot_counter);
    unsigned byte vector_source(snapshot_counter);
    double q0(snapshot_counter);
    double q1(snapshot_counter);
    double q2(snapshot_counter);
    double q3(snapshot_counter);
    double tec(snapshot_counter);
    double geomag_f(snapshot_counter);
    double geomag_d(snapshot_counter);
    double geomag_i(snapshot_counter);
    float sun_ra(snapshot_counter);
    float sun_dec(snapshot_counter);
    float sun_bt(snapshot_counter);
    float accuracy(snapshot_counter);
    float radiometric_accuracy(snapshot_counter, radiometric_accuracy_counter);
    unsigned byte x_band(snapshot_counter);
    unsigned byte software_error_flag(snapshot_counter);
    unsigned byte instrument_error_flag(snapshot_counter);
    unsigned byte adf_error_flag(snapshot_counter);
    unsigned byte calibration_error_flag(snapshot_counter);

// global attributes:
        :title = “TBD ;
        :institution = “TBD ;
        :contact = “TBD” ;
        :creation_date = "Tue Mar 18 11:35:05 UTC 2014" ;
        :total_number_of_grid_points = 2645 ;
}
